library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity processor is 
    port();
end entity processor;

architecture behavioral of processor is

    signal 

begin

end behavioral ; -- behavioral