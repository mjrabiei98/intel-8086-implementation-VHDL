library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;


entity datapath is 
    port ();
end entity datapath;

architecture bwhavioral of datapath is

    -- signal 

begin

end bwhavioral ; -- bwhavioralsab